** Profile: "SCHEMATIC1-AC"  [ D:\DEVELOPWORKSPACE\GITHUB\AudioProject\KC_Amp\KC_BaseBoard\Pspice\KCBaseBoard-PSpiceFiles\SCHEMATIC1\AC.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\DevelopProgramFiles\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 1 50K
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
